//File name=Module name=JTAG_spw  2005-1-18      btltz@mail.china.com      btltz from CASIC,China 
//Description:   JTAG organization for SpaceWire node device ,  Approximate area:
//Origin:        SpaceWire Std - Draft-1 of ESTEC,ESA
//--     TODO:
////////////////////////////////////////////////////////////////////////////////////

/*synthesis translate off*/
`timescale 1ns/10ps
/*synthesis translate on */
module JTAG_spw #()
               ( output TDO,
                 input TDI,
					  input TCK
                );

endmodule